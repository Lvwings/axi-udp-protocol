`timescale 1ns / 1ps
/* -----------------------------------------------------------------------------
 Copyright (c) 2014-2022 All rights reserved
 -----------------------------------------------------------------------------
 Author     : lwings    https://github.com/Lvwings
 File       : lca_4bit.sv
 Create     : 2022-06-22 16:07:04
 Revise     : 2022-06-22 16:07:04
 Language   : Verilog 2001
 -----------------------------------------------------------------------------*/

    module lca_4bit (
        input   [3:0]   a,
        input   [3:0]   b,
        input           cin,
        output  [3:0]   sum,
        output          cout
    );

/*------------------------------------------------------------------------------
--  1-bit Full Adder

    sum     =   a ^ b ^ cin
    cout    =   a & b + cin & (a ^ b)

    Lookahead Carry Adder
    
    sum(i)  =   p(i) ^ c(i)             i = 1...n
    c(i)    =   g(i) + c(i-1) & p(i)    i = 1...n
    c(0)    =   cin
    cout    =   c(n)

    p(i)    =   a(i) ^ b(i)
    g(i)    =   a(i) & b(i)
------------------------------------------------------------------------------*/  

/*------------------------------------------------------------------------------
--  generate p and g
------------------------------------------------------------------------------*/
    logic   [3:0]   p;
    logic   [3:0]   g;

    genvar i;
    generate
        for (i = 0; i < 4; i = i+1) begin
           assign p[i]    =   a[i] ^ b[i];
           assign g[i]    =   a[i] & b[i];   
        end
    endgenerate

/*------------------------------------------------------------------------------
--  generate carry
------------------------------------------------------------------------------*/
    logic   [4:0]   c;

    assign c[1] = g[0] + ( c[0] & p[0] );
    assign c[2] = g[1] + ( (g[0] + ( c[0] & p[0]) ) & p[1] );
    assign c[3] = g[2] + ( (g[1] + ( (g[0] + (c[0] & p[0]) ) & p[1])) & p[2] );
    assign c[4] = g[3] + ( (g[2] + ( (g[1] + ( (g[0] + (c[0] & p[0]) ) & p[1])) & p[2] )) & p[3]);
    
    assign c[0] = cin;
    assign cout = c[4];

/*------------------------------------------------------------------------------
--  generate sum 
------------------------------------------------------------------------------*/
     generate
        for (i = 0; i < 4; i = i+1) begin
           assign sum[i]    =   p[i] ^ c[i]; 
        end
    endgenerate   

endmodule : lca_4bit
